/home/jay/openrisc/minsoc/prj/../rtl/verilog/adv_debug_sys/Hardware/altera_virtual_jtag/rtl/vhdl//altera_virtual_jtag.vhd
